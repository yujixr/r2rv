parameter RAM_SIZE_LOG = 8;
parameter RAM_SIZE = 2**RAM_SIZE_LOG;

module writer(
  input logic clk,
  input logic [31:0] RAM_READ[RAM_SIZE-1:0],
  output logic [31:0] RAM_WRITE[RAM_SIZE-1:0],
  input logic enabler,
  input ldst_mode mode,
  input logic [RAM_SIZE_LOG-1:0] addr,
  input logic [31:0] data
);

genvar i;
generate
  for (i = 0; i < RAM_SIZE; i++) begin: Update
    always_ff @(negedge clk)
      if ((addr==i) & enabler)
        RAM_WRITE[i] <= data;
      else
        RAM_WRITE[i] <= RAM_READ[i];
  end
endgenerate

endmodule


module reader(
  input logic [31:0] RAM[RAM_SIZE-1:0],
  input ldst_mode mode,
  input logic [RAM_SIZE_LOG-1:0] addr,
  output logic [31:0] data
);

assign data = RAM[addr];

endmodule


module mem(
  input logic clk, we,
  input logic [31:0] ra1, ra2, wa3,
  input ldst_mode rm1, rm2, wm3,
  input logic [31:0] wd3,
  output logic [31:0] rd1, rd2,
  output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5
);

logic [31:0] imem[RAM_SIZE-1:0], dmem[RAM_SIZE-1:0], stdout;

initial begin
  $readmemh("imem.dat", imem);
  $readmemh("dmem.dat", dmem);
end

reader read1(imem, rm1, ra1[RAM_SIZE_LOG+1:2], rd1);
reader read2(dmem, rm2, ra2[RAM_SIZE_LOG+1:2], rd2);
writer write(clk, dmem, dmem, we, wm3, wa3[RAM_SIZE_LOG+1:2], wd3);

assign stdout = dmem['h3f];

hex_display hex2023(stdout[23:20], HEX5);
hex_display hex1619(stdout[19:16], HEX4);
hex_display hex1215(stdout[15:12], HEX3);
hex_display hex0811(stdout[11:8], HEX2);
hex_display hex0407(stdout[7:4], HEX1);
hex_display hex0003(stdout[3:0], HEX0);

endmodule
